module RandomGenerator (
        input wire clk,
        input wire reset,
        input [15:0] seed,
        output [15:0] random_number
    );
    reg [15:0] lfsr;

    always @(posedge clk or posedge reset) begin
        if (reset) begin
            lfsr <= seed;
        end
        else begin
            lfsr <= {lfsr[14:0], lfsr[15] ^ lfsr[14]};
        end
    end

    assign random_number = lfsr;
endmodule
